`timescale 1ns / 1ps

/// \brief Template interface for VeSPA Custom Bus slave device
/// \input i_Clk Source Clock signal for the slave device, logic is processed on rising edges of this signal
/// \input i_Rst Reset signal for the device, active high
/// \input i_WEnable Write Enable signal. If this signal is set to high during a rising edge of the clock,
/// data is writen to the slave register file
/// \input i_WAddr Address of the register file that data should be writen to. This is a virtual address,
/// that should be generated by a Bus Interconnect device
/// \input i_WData Data writen to the slave register file if all the required conditions are complied
/// \input i_REnable Read Enable signal. If this signal is set to high during a rising edge of the clock,
/// data is read from the slave register file
/// \input i_RAddr Address of the register file that data will be read from. Simmilar to the i_WAddr, this
/// address should be generated by a Bus Interconnect device
/// \output o_RData When a read operation occurs, data is put on this output
/// \output o_Err This signal indicated an internal error occured on the device, such as an invalid address
module SlaveInterface
(
    //Bus related signals
    input i_Clk,
    input i_Rst,
    input i_WEnable,
    input [31:0] i_WAddr,
    input [31:0] i_WData,
    input i_REnable,
    input [31:0] i_RAddr,
    output [31:0] o_RData,
    output reg o_Err,
    //User signals begin here
    output o_MemBusy
);

wire [31:0] w_MemAddr;
wire [3:0] w_WEnA;
wire w_RstA, w_RstB;

assign w_MemAddr = i_WEnable ? i_WAddr : i_REnable ? i_RAddr : 0;
assign w_WEnA = {i_WEnable, i_WEnable, i_WEnable, i_WEnable};

VeSPA_RAM _Bram(
  .clka(i_Clk),
  .rsta(i_Rst),
  .wea(w_WEnA),
  .addra(w_MemAddr),
  .dina(i_WData),
  .douta(o_RData),
  .rsta_busy(o_MemBusy)
);

endmodule
